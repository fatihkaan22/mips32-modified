module shift_left_2(a, o);
input [31:0] a;
output [31:0] o;

buf b0(o[0],1'b0),
    b1(o[1], 1'b0),
    b2(o[2], a[0]),
    b3(o[3], a[1]),
    b4(o[4], a[2]),
    b5(o[5], a[3]),
    b6(o[6], a[4]),
    b7(o[7], a[5]),
    b8(o[8], a[6]),
    b9(o[9], a[7]),
    b10(o[10], a[8]),
    b11(o[11], a[9]),
    b12(o[12], a[10]),
    b13(o[13], a[11]),
    b14(o[14], a[12]),
    b15(o[15], a[13]),
    b16(o[16], a[14]),
    b17(o[17], a[15]),
    b18(o[18], a[16]),
    b19(o[19], a[17]),
    b20(o[20], a[18]),
    b21(o[21], a[19]),
    b22(o[22], a[20]),
    b23(o[23], a[21]),
    b24(o[24], a[22]),
    b25(o[25], a[23]),
    b26(o[26], a[24]),
    b27(o[27], a[25]),
    b28(o[28], a[26]),
    b29(o[29], a[27]),
    b30(o[30], a[28]),
    b31(o[31], a[29]);

endmodule
